library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity cordic_postprocess is
    port (
        clk   : in std_logic;
        reset : in std_logic

    );
end entity cordic_postprocess;

architecture rtl of cordic_postprocess is

begin

end architecture;